module mux(
    
);

endmodule