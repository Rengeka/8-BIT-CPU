module decoder(
    
);

endmodule